library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity useVcc is
    port (
    output : out std_logic

    );
end useVcc;

architecture structural of useVcc is



begin
     output <= '1';
end structural;